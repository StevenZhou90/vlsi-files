magic
tech scmos
timestamp 1759278974
<< error_p >>
rect 121 306 440 404
rect 121 4 440 57
<< metal1 >>
rect 12 1289 13 1294
rect 18 1289 42 1294
rect 33 1102 35 1107
rect 12 1012 13 1017
rect 18 1012 43 1017
rect 12 915 13 920
rect 18 915 42 920
rect 12 638 13 643
rect 18 638 43 643
rect 18 541 40 546
rect 17 264 40 269
<< m123contact >>
rect 37 1476 42 1481
rect 13 1289 18 1294
rect 35 1199 40 1204
rect 35 1102 40 1107
rect 13 1012 18 1017
rect 13 915 18 920
rect 35 825 40 830
rect 37 728 42 733
rect 13 638 18 643
rect 12 541 18 546
rect 36 451 42 456
rect 33 352 40 359
rect 12 264 17 269
rect 33 77 40 84
<< metal3 >>
rect 33 1476 37 1481
rect 12 1289 13 1294
rect 12 1017 18 1289
rect 33 1204 40 1476
rect 33 1199 35 1204
rect 12 1012 13 1017
rect 33 1102 35 1107
rect 12 915 13 920
rect 12 643 18 915
rect 33 830 40 1102
rect 33 825 35 830
rect 12 638 13 643
rect 33 728 37 733
rect 12 269 18 541
rect 33 456 40 728
rect 33 451 36 456
rect 17 264 18 269
rect 33 84 40 352
use shift  shift_0
timestamp 1759278974
transform 1 0 40 0 1 4
box -36 0 400 1477
<< end >>
