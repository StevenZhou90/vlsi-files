magic
tech scmos
timestamp 1758948824
use fblock_one  fblock_one_0
array 0 7 173 0 0 227
timestamp 1758948824
transform 1 0 -15 0 1 28
box 15 -28 177 201
<< end >>
