magic
tech scmos
timestamp 1758765833
<< error_s >>
rect 68 -44 72 -43
rect 65 -46 72 -44
rect 62 -47 72 -46
rect 63 -51 68 -47
<< metal1 >>
rect 72 163 77 181
rect 40 146 54 152
rect 40 136 47 146
rect 68 144 77 149
rect 89 146 101 152
rect 32 124 40 129
rect 68 113 73 144
rect 94 138 101 146
rect 30 98 35 106
rect 51 89 57 96
rect 51 70 56 89
rect 33 65 56 70
rect 85 70 90 95
rect 95 84 102 89
rect 107 84 108 89
rect 85 65 109 70
rect 5 50 12 54
rect 33 41 38 65
rect 16 10 22 26
rect 50 24 55 29
rect 5 -7 12 8
rect 49 13 55 23
rect 49 8 50 13
rect 87 15 93 23
rect 104 22 109 65
rect 112 60 117 74
rect 130 65 136 89
rect 130 57 137 65
rect 131 48 136 57
rect 92 10 93 15
rect 49 4 55 8
rect 120 9 126 24
rect 26 1 30 4
rect 96 1 101 6
rect 26 -4 101 1
rect -17 -12 158 -7
rect -1 -35 8 -30
rect 39 -35 46 -30
rect 93 -35 104 -30
rect 129 -35 142 -30
rect -17 -51 62 -47
rect 68 -51 158 -47
rect -17 -52 158 -51
rect -6 -63 -1 -60
rect 34 -63 39 -60
rect 104 -63 109 -60
rect 142 -63 147 -60
<< m2contact >>
rect 40 125 47 130
rect 120 125 125 130
rect 13 102 18 107
rect 76 102 81 107
rect 114 101 119 106
rect 131 101 136 106
rect 30 93 35 98
rect 60 93 65 98
rect 19 84 24 89
rect 102 84 107 89
rect 112 74 117 79
rect 5 54 12 61
rect 96 52 101 57
rect 60 43 65 48
rect 6 28 11 33
rect 77 28 82 33
rect 16 4 22 10
rect 41 4 46 9
rect 131 43 136 48
rect 112 4 117 9
rect 121 4 127 9
rect -6 -35 -1 -30
rect 20 -35 25 -30
rect 34 -35 39 -30
rect 104 -35 109 -30
rect 116 -35 121 -30
rect 142 -35 147 -30
rect -6 -60 -1 -55
rect 34 -60 39 -55
rect 104 -60 109 -55
rect 142 -60 147 -55
<< metal2 >>
rect 1 125 40 130
rect 47 125 120 130
rect 1 76 8 125
rect 18 102 76 107
rect 35 93 60 98
rect 24 84 102 89
rect 114 79 119 101
rect 1 69 12 76
rect 117 74 119 79
rect 5 61 12 69
rect 131 57 136 101
rect 101 52 136 57
rect 65 43 131 48
rect 11 28 77 33
rect 16 -13 22 4
rect 41 1 46 4
rect 112 1 117 4
rect 41 -4 117 1
rect 121 -8 127 4
rect 16 -19 25 -13
rect 20 -30 25 -19
rect 116 -14 127 -8
rect 116 -30 121 -14
rect -6 -55 -1 -35
rect 34 -55 39 -35
rect 104 -55 109 -35
rect 142 -55 147 -35
<< m123contact >>
rect 50 8 55 13
rect 87 10 92 15
rect 60 5 65 10
rect 58 -35 63 -30
rect 79 -35 84 -30
rect 62 -51 68 -47
<< metal3 >>
rect 50 1 55 8
rect 65 5 74 10
rect 50 -4 63 1
rect 58 -30 63 -4
rect 68 -47 74 5
rect 87 1 92 10
rect 79 -4 92 1
rect 79 -30 84 -4
use inv  inv_3
timestamp 1758764680
transform -1 0 129 0 1 -48
box -9 -7 21 44
use inv  inv_0
timestamp 1758764680
transform 1 0 12 0 1 -48
box -9 -7 21 44
use inv  inv_1
timestamp 1758764680
transform 1 0 50 0 1 -48
box -9 -7 21 44
use inv  inv_2
timestamp 1758764680
transform -1 0 92 0 1 -48
box -9 -7 21 44
use tgmux2  tgmux2_0
timestamp 1758764680
transform 1 0 20 0 1 16
box -20 -16 51 47
use tgmux2  tgmux2_1
timestamp 1758764680
transform 1 0 91 0 1 16
box -20 -16 51 47
use inv  inv_5
timestamp 1758764680
transform -1 0 127 0 1 88
box -9 -7 21 44
use inv  inv_4
timestamp 1758764680
transform -1 0 26 0 1 88
box -9 -7 21 44
use tgmux2  tgmux2_2
timestamp 1758764680
transform 1 0 55 0 1 93
box -20 -16 51 47
use inv  inv_6
timestamp 1758764680
transform 0 -1 90 1 0 155
box -9 -7 21 44
<< labels >>
rlabel metal1 42 144 42 144 1 Vdd!
rlabel metal1 95 143 95 143 1 GND!
rlabel metal1 73 179 73 179 5 f
rlabel metal2 37 95 37 95 1 a
rlabel metal2 133 94 133 94 1 b
rlabel metal2 37 105 37 105 1 bara
rlabel metal2 116 81 116 81 1 barb
rlabel metal1 35 -62 35 -62 1 g1
rlabel metal1 106 -62 106 -62 1 g2
rlabel metal1 96 67 96 67 1 t1
rlabel metal1 43 68 43 68 1 t0
rlabel metal1 -5 -62 -5 -62 1 g0
rlabel metal1 143 -62 143 -62 1 g3
rlabel metal1 128 -49 128 -49 5 Vdd!
rlabel metal1 13 -49 13 -49 5 Vdd!
rlabel metal1 51 -49 51 -49 5 Vdd!
rlabel metal1 91 -49 91 -49 5 Vdd!
<< end >>
