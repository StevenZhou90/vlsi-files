magic
tech scmos
timestamp 1759201369
<< metal1 >>
rect -20 129 121 134
rect 251 99 261 104
rect -19 93 121 98
rect -19 73 -14 78
rect 106 64 167 69
rect 106 52 111 64
rect 121 48 126 61
rect 111 43 126 48
rect -19 37 -14 42
rect 207 12 212 59
rect 106 7 212 12
rect -19 0 -14 5
use mux2  mux2_1
timestamp 1759197544
transform -1 0 382 0 -1 130
box 126 -4 261 74
use mux2  mux2_0
timestamp 1759197544
transform -1 0 242 0 -1 74
box 126 -4 261 74
<< labels >>
rlabel metal1 -17 39 -17 39 3 u
rlabel metal1 -17 3 -17 3 2 au
rlabel metal1 -16 76 -16 76 3 ad
rlabel metal1 -17 95 -17 95 3 s
rlabel metal1 -18 132 -18 132 4 a
rlabel metal1 258 101 258 101 7 out
<< end >>
