magic
tech scmos
timestamp 1759374011
<< metal1 >>
rect 137 215 144 220
rect 137 208 149 215
rect 558 208 565 220
rect 979 208 986 220
rect 1400 208 1407 220
rect 1821 208 1828 220
rect 2242 208 2249 220
rect 2663 208 2670 220
rect 3084 208 3091 220
rect 187 149 192 169
rect 608 149 613 169
rect 1029 149 1034 169
rect 1450 149 1455 169
rect 1871 149 1876 169
rect 2292 149 2297 169
rect 2713 149 2718 169
rect 3134 149 3139 169
rect 7 140 15 143
rect 368 92 413 96
rect 7 -1 15 2
<< metal2 >>
rect -12 188 -7 247
rect 0 204 5 247
rect -1 199 18 204
rect 52 194 57 199
rect 409 188 414 247
rect 421 204 426 247
rect 421 199 439 204
rect 830 188 835 247
rect 842 204 847 247
rect 842 199 860 204
rect 1251 188 1256 247
rect 1263 204 1268 247
rect 1263 199 1281 204
rect 1672 188 1677 247
rect 1684 204 1689 247
rect 1684 199 1702 204
rect 2093 188 2098 247
rect 2105 204 2110 247
rect 2105 199 2123 204
rect 2514 188 2519 247
rect 2526 204 2531 247
rect 2526 199 2544 204
rect 2935 188 2940 247
rect 2947 204 2952 247
rect 2947 199 2965 204
rect -12 183 5 188
rect 409 183 426 188
rect 830 183 847 188
rect 1251 183 1268 188
rect 1672 183 1689 188
rect 2093 183 2110 188
rect 2514 183 2531 188
rect 2935 183 2952 188
rect 0 110 5 183
rect 421 111 426 183
rect 0 107 9 110
rect 0 106 5 107
rect 421 106 447 111
rect 842 111 847 183
rect 842 106 888 111
rect 1263 111 1268 183
rect 1263 106 1309 111
rect 1684 111 1689 183
rect 1684 106 1730 111
rect 2105 111 2110 183
rect 2105 106 2151 111
rect 2526 111 2531 183
rect 2526 106 2572 111
rect 2947 111 2952 183
rect 2947 106 2993 111
rect 0 12 26 18
rect 3230 17 3368 23
<< m123contact >>
rect 171 225 176 230
rect 144 215 149 220
rect 52 199 57 204
rect 592 225 597 230
rect 565 215 570 220
rect 473 199 478 204
rect 1013 225 1018 230
rect 986 215 991 220
rect 894 199 899 204
rect 1434 225 1439 230
rect 1407 215 1412 220
rect 1315 199 1320 204
rect 1855 225 1860 230
rect 1828 215 1833 220
rect 1736 199 1741 204
rect 2276 225 2281 230
rect 2249 215 2254 220
rect 2157 199 2162 204
rect 2697 225 2702 230
rect 2670 215 2675 220
rect 2578 199 2583 204
rect 3118 225 3123 230
rect 3091 215 3096 220
rect 2999 199 3004 204
rect 385 110 390 115
rect 806 110 811 115
rect 1227 110 1232 115
rect 1648 110 1653 115
rect 2069 110 2074 115
rect 2490 110 2495 115
rect 2911 110 2916 115
rect 3332 110 3337 115
<< metal3 >>
rect 52 234 3004 239
rect 52 204 57 234
rect 51 199 52 204
rect 51 153 57 199
rect 144 160 149 215
rect 26 147 57 153
rect 74 155 149 160
rect 74 148 79 155
rect 171 148 176 225
rect 473 204 478 234
rect 565 160 570 215
rect 495 155 570 160
rect 592 148 597 225
rect 894 204 899 234
rect 986 160 991 215
rect 916 155 991 160
rect 1013 148 1018 225
rect 1315 204 1320 234
rect 1407 160 1412 215
rect 1337 155 1412 160
rect 1434 148 1439 225
rect 1736 204 1741 234
rect 1828 160 1833 215
rect 1758 155 1833 160
rect 1855 148 1860 225
rect 2157 204 2162 234
rect 2249 160 2254 215
rect 2179 155 2254 160
rect 2276 148 2281 225
rect 2578 204 2583 234
rect 2670 160 2675 215
rect 2600 155 2675 160
rect 2697 148 2702 225
rect 2999 204 3004 234
rect 3091 160 3096 215
rect 3021 155 3096 160
rect 3118 148 3123 225
rect 26 12 32 147
rect 385 -17 390 110
rect 806 -17 811 110
rect 1227 -17 1232 110
rect 1648 -17 1653 110
rect 2069 -17 2074 110
rect 2490 -17 2495 110
rect 2911 -17 2916 110
rect 3332 -17 3337 110
use xor3  xor3_0
array 0 7 421 0 0 -70
timestamp 1759372879
transform 1 0 95 0 -1 171
box -95 -76 100 16
use addsub_one  addsub_one_0
array 0 7 421 0 0 158
timestamp 1759372879
transform 1 0 28 0 1 63
box -28 -66 393 92
<< labels >>
rlabel metal2 425 200 425 200 1 b1
rlabel metal2 845 201 845 201 1 b2
rlabel metal2 1266 201 1266 201 1 b3
rlabel metal2 1686 201 1686 201 1 b4
rlabel metal2 2108 201 2108 201 1 b5
rlabel metal2 2530 202 2530 202 1 b6
rlabel metal2 2951 201 2951 201 1 b7
rlabel metal1 9 141 9 141 1 Vdd!
rlabel metal1 10 1 10 1 1 GND!
rlabel metal2 845 108 845 108 1 a2
rlabel metal2 1264 108 1264 108 1 a3
rlabel metal2 1686 108 1686 108 1 a4
rlabel metal2 2108 108 2108 108 1 a5
rlabel metal2 2531 108 2531 108 1 a6
rlabel metal2 2951 108 2951 108 1 a7
rlabel metal2 3355 20 3355 20 1 cout
rlabel metal2 3 14 3 14 3 cin
rlabel metal2 5 201 5 201 3 b0
rlabel metal2 426 201 426 201 3 b1
rlabel metal2 847 201 847 201 3 b2
rlabel metal2 1268 201 1268 201 3 b3
rlabel metal2 1689 201 1689 201 3 b4
rlabel metal2 2110 201 2110 201 3 b5
rlabel metal2 2531 201 2531 201 3 b6
rlabel metal2 2952 201 2952 201 3 b7
rlabel metal2 4 109 4 109 3 a0
rlabel metal2 425 109 425 109 3 a1
rlabel metal2 846 109 846 109 3 a2
rlabel metal2 1267 109 1267 109 3 a3
rlabel metal2 1688 109 1688 109 3 a4
rlabel metal2 2109 109 2109 109 3 a5
rlabel metal2 2530 109 2530 109 3 a6
rlabel metal2 2951 109 2951 109 3 a7
rlabel metal3 386 -15 386 -15 1 s0
rlabel metal3 807 -15 807 -15 1 s1
rlabel metal3 1228 -15 1228 -15 1 s2
rlabel metal3 1650 -14 1650 -14 1 s3
rlabel metal3 2070 -15 2070 -15 1 s4
rlabel metal3 2491 -14 2491 -14 1 s5
rlabel metal3 2912 -14 2912 -14 1 s6
rlabel metal3 3334 -14 3334 -14 1 s7
<< end >>
