magic
tech scmos
timestamp 1758735917
<< nwell >>
rect -9 16 21 44
<< pwell >>
rect -9 -7 21 16
<< ntransistor >>
rect 5 5 7 10
<< ptransistor >>
rect 5 22 7 32
<< ndiffusion >>
rect 4 5 5 10
rect 7 5 8 10
<< pdiffusion >>
rect 3 22 5 32
rect 7 22 8 32
<< ndcontact >>
rect -1 5 4 10
rect 8 5 13 10
<< pdcontact >>
rect -2 22 3 32
rect 8 22 13 32
<< psubstratepcontact >>
rect -6 -4 -1 1
rect 13 -4 18 1
<< nsubstratencontact >>
rect -6 36 -1 41
rect 13 36 18 41
<< polysilicon >>
rect 5 32 7 35
rect 5 15 7 22
rect 5 2 7 5
<< polycontact >>
rect 0 13 5 18
<< polynplus >>
rect 5 10 7 15
<< metal1 >>
rect -9 36 -6 41
rect -1 36 13 41
rect 18 36 21 41
rect -2 32 3 36
rect -9 13 0 18
rect 8 10 13 22
rect -1 1 4 5
rect -9 -4 -6 1
rect -1 -4 13 1
rect 18 -4 21 1
<< labels >>
rlabel metal1 -7 14 -7 14 3 in
rlabel metal1 9 15 9 15 1 out
rlabel metal1 1 39 1 39 5 Vdd!
rlabel metal1 2 -3 2 -3 1 GND!
<< end >>
