magic
tech scmos
timestamp 1759005747
<< metal1 >>
rect 231 69 261 74
rect 166 62 174 67
rect 205 62 211 67
rect 156 51 161 58
rect 170 30 175 43
rect 215 30 220 43
rect 249 37 254 38
rect 231 29 236 34
rect 249 32 261 37
rect 249 29 254 32
rect 220 12 226 17
rect 197 1 202 2
rect 231 -4 261 1
<< m2contact >>
rect 192 69 197 74
rect 226 69 231 74
rect 200 60 205 65
rect 161 51 166 56
rect 235 52 240 57
rect 162 40 167 45
rect 131 35 136 40
rect 146 35 151 40
rect 126 26 131 31
rect 197 38 202 43
rect 192 29 197 34
rect 249 38 254 43
rect 226 29 231 34
rect 146 17 151 22
rect 200 20 205 25
rect 215 12 220 17
rect 197 -4 202 1
rect 226 -4 231 1
<< metal2 >>
rect 197 69 226 74
rect 131 60 200 65
rect 131 40 136 60
rect 166 52 235 56
rect 166 51 240 52
rect 146 31 151 35
rect 131 26 151 31
rect 162 25 167 40
rect 202 38 249 43
rect 197 29 226 34
rect 162 20 200 25
rect 146 11 151 17
rect 215 11 220 12
rect 146 6 220 11
rect 202 -4 226 1
use nand2  nand2_1
timestamp 1759005747
transform 0 -1 221 1 0 3
box -7 -2 29 54
use nand2  nand2_0
timestamp 1759005747
transform 0 -1 221 1 0 45
box -7 -2 29 54
use nand2  nand2_2
timestamp 1759005747
transform 1 0 138 0 1 16
box -7 -2 29 54
use inv  inv_0
timestamp 1759005747
transform -1 0 244 0 1 16
box -9 -7 21 44
<< labels >>
rlabel space 217 59 217 59 1 GND!
rlabel metal1 172 36 172 36 1 Vdd!
rlabel metal1 257 -2 257 -2 8 A
rlabel metal1 257 71 257 71 6 B
rlabel metal1 258 34 258 34 7 SEL
rlabel m2contact 127 28 127 28 3 OUT
<< end >>
