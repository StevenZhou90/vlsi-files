magic
tech scmos
timestamp 1759289494
<< metal1 >>
rect 0 1473 6 1500
rect -45 1436 7 1441
rect -45 1254 -40 1436
rect 0 1286 6 1313
rect 42 1290 47 1315
rect 87 1290 92 1315
rect -45 1249 8 1254
rect -45 1067 -40 1249
rect 0 1099 6 1126
rect 42 1102 47 1127
rect 87 1103 92 1128
rect -45 1062 6 1067
rect -45 880 -40 1062
rect 0 912 6 939
rect 42 916 47 941
rect 87 916 92 941
rect -45 875 6 880
rect -45 693 -40 875
rect 0 725 6 752
rect 42 729 47 754
rect 87 729 92 754
rect -45 688 6 693
rect -45 506 -40 688
rect 0 538 6 565
rect 42 542 47 567
rect 87 542 92 567
rect -45 501 6 506
rect -45 319 -40 501
rect 0 355 6 378
rect 42 355 47 380
rect 87 355 92 380
rect 0 351 1 355
rect -45 314 6 319
rect -45 132 -40 314
rect 0 164 6 191
rect 42 168 47 193
rect 87 168 92 193
rect -45 127 6 132
rect 5 73 16 78
<< metal2 >>
rect -35 1340 16 1345
rect -35 1158 -30 1340
rect -35 1153 16 1158
rect -35 971 -30 1153
rect -35 966 16 971
rect -35 784 -30 966
rect -35 779 16 784
rect -35 597 -30 779
rect -35 592 16 597
rect -35 410 -30 592
rect -35 405 16 410
rect -35 223 -30 405
rect -35 218 16 223
rect -35 36 -30 218
rect -35 31 16 36
<< m123contact >>
rect 1 350 6 355
rect 0 73 5 78
<< metal3 >>
rect -17 1008 -12 1290
rect 18 1195 23 1477
rect -17 634 -12 916
rect 18 821 23 1103
rect -17 260 -12 542
rect 18 447 23 729
rect 0 350 1 355
rect 6 350 23 355
rect 18 78 23 350
rect 5 73 23 78
use shift_one  shift_one_0
array 0 0 144 0 7 187
timestamp 1759289462
transform 1 0 -2 0 1 7
box 2 -7 146 161
<< end >>
