magic
tech scmos
timestamp 1758767863
<< nwell >>
rect -7 24 29 54
<< pwell >>
rect -7 -2 29 24
<< ntransistor >>
rect 5 10 7 16
rect 14 10 16 16
<< ptransistor >>
rect 5 30 7 42
rect 14 30 16 42
<< ndiffusion >>
rect 4 10 5 16
rect 7 10 14 16
rect 16 10 17 16
<< pdiffusion >>
rect 4 35 5 42
rect -1 30 5 35
rect 7 35 14 42
rect 7 30 8 35
rect 13 30 14 35
rect 16 35 18 42
rect 16 30 23 35
<< ndcontact >>
rect -1 10 4 16
rect 17 10 22 16
<< pdcontact >>
rect -1 35 4 42
rect 8 30 13 35
rect 18 35 23 42
<< psubstratepcontact >>
rect 0 1 5 6
rect 18 1 23 6
<< nsubstratencontact >>
rect 2 46 7 51
rect 16 46 21 51
<< polysilicon >>
rect 5 42 7 45
rect 14 42 16 45
rect 5 16 7 30
rect 14 16 16 30
rect 5 7 7 10
rect 14 7 16 10
<< polycontact >>
rect 0 19 5 24
rect 16 24 21 29
<< metal1 >>
rect -7 46 2 51
rect 7 46 16 51
rect 21 46 29 51
rect -1 42 4 46
rect 18 42 23 46
rect -7 19 0 24
rect 8 21 13 30
rect 21 24 29 29
rect 8 17 22 21
rect 17 16 22 17
rect -1 6 4 10
rect -7 1 0 6
rect 5 1 18 6
rect 23 1 29 6
<< labels >>
rlabel metal1 -1 49 -1 49 4 Vdd!
rlabel metal1 20 18 20 18 1 out
rlabel metal1 -1 2 -1 2 2 GND!
rlabel metal1 -5 20 -5 20 3 A
rlabel metal1 23 25 23 25 7 B
<< end >>
