magic
tech scmos
timestamp 1759364525
<< metal1 >>
rect -27 77 80 82
rect 189 77 203 82
rect 363 77 393 82
rect 198 71 203 77
rect 13 66 14 71
rect 198 66 209 71
rect 141 41 149 45
rect 145 31 149 41
rect 187 43 192 48
rect 197 43 199 48
rect 333 45 337 50
rect 187 31 191 43
rect 333 41 344 45
rect 333 39 337 41
rect 340 33 344 41
rect 145 27 191 31
rect 198 26 209 31
rect 340 29 385 33
rect 198 22 203 26
rect -1 17 80 21
rect 190 17 203 22
rect -1 -60 3 17
rect 101 -9 128 -4
rect 157 -9 198 -4
rect 195 -16 198 -9
rect 99 -39 101 -34
rect 157 -38 192 -34
rect 157 -39 198 -38
rect 189 -43 198 -39
rect 227 -45 250 -41
rect 101 -54 128 -49
rect 70 -60 75 -54
rect -27 -64 75 -60
rect 159 -61 164 -49
rect 233 -59 238 -56
rect 159 -66 202 -61
rect 233 -64 393 -59
<< m2contact >>
rect 192 43 197 48
rect 199 43 204 48
rect 159 -31 164 -26
rect 70 -36 75 -31
rect 128 -36 133 -31
rect 250 -46 255 -41
<< metal2 >>
rect -27 43 12 48
rect 7 -31 12 43
rect 192 39 197 43
rect 192 12 196 39
rect 118 8 196 12
rect 7 -36 70 -31
rect 118 -32 122 8
rect 164 -1 242 4
rect 164 -2 247 -1
rect 164 -31 170 -2
rect 118 -36 128 -32
rect 159 -32 170 -31
rect 164 -45 170 -32
rect 254 -41 393 -40
rect -27 -51 170 -45
rect 255 -46 393 -41
rect 387 -51 393 -46
<< m3contact >>
rect 47 43 52 48
rect 242 43 247 48
rect 242 -1 247 4
<< m123contact >>
rect 8 66 13 71
rect 70 -9 75 -4
rect 101 -28 106 -23
rect 101 -39 106 -34
rect 229 -38 234 -33
<< metal3 >>
rect 8 -4 13 66
rect 46 43 47 48
rect 46 17 52 43
rect 22 11 52 17
rect 39 6 45 11
rect 39 0 114 6
rect 8 -9 70 -4
rect 108 -23 114 0
rect 242 4 247 43
rect 106 -28 114 -23
rect 106 -58 111 -34
rect 234 -38 245 -33
rect 240 -58 245 -38
rect 106 -63 245 -58
use nand2  nand2_2
timestamp 1759005747
transform 1 0 205 0 1 -62
box -7 -2 29 54
use nand2  nand2_1
timestamp 1759005747
transform 1 0 135 0 1 -55
box -7 -2 29 54
use nand2  nand2_0
timestamp 1759005747
transform 1 0 77 0 1 -55
box -7 -2 29 54
use xor3  xor3_1
timestamp 1759285841
transform 1 0 290 0 1 76
box -95 -76 100 16
use xor3  xor3_0
timestamp 1759285841
transform 1 0 95 0 1 76
box -95 -76 100 16
<< labels >>
rlabel metal2 -27 43 12 48 1 a
rlabel metal3 39 0 114 6 1 b
rlabel metal2 -27 -51 170 -45 1 cin
rlabel metal2 255 -46 393 -40 1 cout
rlabel metal1 340 29 385 33 1 s
<< end >>
