magic
tech scmos
timestamp 1759286262
<< error_p >>
rect 117 302 436 400
rect 117 0 436 53
use shift2  shift2_0
timestamp 1759286262
transform 1 0 -4 0 1 -4
box 4 4 440 1481
<< end >>
