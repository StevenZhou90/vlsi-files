magic
tech scmos
timestamp 1759005747
<< metal1 >>
rect 156 159 164 164
rect 25 153 34 158
rect 36 106 41 149
rect 73 123 78 128
rect 73 118 86 123
rect 81 107 86 118
rect 91 68 101 73
rect 90 23 100 28
rect 15 -28 20 -18
rect 88 -28 93 -18
rect 99 -28 104 -18
rect 172 -28 177 -18
<< metal2 >>
rect 129 123 134 128
rect 57 -11 146 -6
<< m123contact >>
rect 129 196 134 201
rect 100 165 105 170
rect 100 123 105 128
rect 45 112 50 117
rect 129 112 134 117
<< metal3 >>
rect 105 165 124 168
rect 100 163 124 165
rect 45 123 100 128
rect 45 117 50 123
rect 119 -18 124 163
rect 129 117 134 196
use mux2  mux2_0
timestamp 1759005747
transform 0 1 19 -1 0 243
box 126 -4 261 74
use mux2  mux2_1
timestamp 1759005747
transform 0 1 103 -1 0 243
box 126 -4 261 74
use mux2  mux2_2
timestamp 1759005747
transform 1 0 -97 0 1 127
box 126 -4 261 74
<< labels >>
rlabel metal1 161 162 161 162 1 A
rlabel metal1 26 155 26 155 1 OUT
rlabel metal1 17 -26 17 -26 2 g0
rlabel metal1 89 -26 89 -26 1 g1
rlabel metal1 100 -26 100 -26 1 g2
rlabel metal1 173 -26 173 -26 8 g3
rlabel metal2 84 -8 84 -8 1 B
<< end >>
