magic
tech scmos
timestamp 1758768781
<< nwell >>
rect -4 29 32 66
<< pwell >>
rect -4 -2 32 29
<< ntransistor >>
rect 9 10 11 22
rect 18 10 20 22
<< ptransistor >>
rect 9 35 11 53
rect 18 35 20 53
<< ndiffusion >>
rect 3 17 9 22
rect 8 10 9 17
rect 11 15 12 22
rect 17 15 18 22
rect 11 10 18 15
rect 20 17 26 22
rect 20 10 21 17
<< pdiffusion >>
rect 7 46 9 53
rect 2 35 9 46
rect 11 35 18 53
rect 20 42 26 53
rect 20 35 21 42
<< ndcontact >>
rect 3 10 8 17
rect 12 15 17 22
rect 21 10 26 17
<< pdcontact >>
rect 2 46 7 53
rect 21 35 26 42
<< psubstratepcontact >>
rect 3 1 8 6
rect 21 1 26 6
<< nsubstratencontact >>
rect 4 57 9 62
rect 17 57 22 62
<< polysilicon >>
rect 9 53 11 56
rect 18 53 20 56
rect 9 22 11 35
rect 18 22 20 35
rect 9 7 11 10
rect 18 7 20 10
<< polycontact >>
rect 4 23 9 28
rect 20 23 25 28
<< metal1 >>
rect -4 57 4 62
rect 9 57 17 62
rect 22 57 32 62
rect 2 53 7 57
rect 12 31 26 35
rect 0 23 4 28
rect 12 22 17 31
rect 25 23 29 28
rect 3 6 8 10
rect 21 6 26 10
rect -2 1 3 6
rect 8 1 21 6
rect 26 1 30 6
<< labels >>
rlabel metal1 11 3 11 3 1 GND!
rlabel nwell 10 60 10 60 5 Vdd!
rlabel metal1 18 34 18 34 1 out
rlabel polycontact 22 25 22 25 1 B
rlabel polycontact 7 25 7 25 1 A
<< end >>
